module InstMem(Addr, Inst, clk, set);
  input[15:0] Addr;
  input clk, set;
  output [15:0] Inst;
  
  reg [15:0] InstMem [0:1024*64-1];
  
  assign Inst = 
			(Addr == 'd0 ) ? 'b1001_001_000_000_101: // addi r1 = 5	
			(Addr == 'd1 ) ? 'b1001_010_000_111_011: // addi r2 = -5	
			(Addr == 'd2 ) ? 'b1001_011_010_001_111: // addi r3 = R2 +15 = 10
			(Addr == 'd3 ) ? 'b1001_100_010_111_111: // addi r4 = R2 - 1 = -6
			(Addr == 'd4 ) ? 'b1001_101_010_000_101: // addi r5 = R2 + 5 = 0
			(Addr == 'd5 ) ? 'b0000_111_100_101_000: //nop
			(Addr == 'd6 ) ? 'b1001_110_101_000_110: // addi r6 = R5 + 6 = 6
			(Addr == 'd7 ) ? 'b0000_000_000_000_000: //nop
			(Addr == 'd8 ) ? 'b0000_000_000_000_000: //nop
			(Addr == 'd9 ) ? 'b1001_111_110_000_101: // addi r7 = R6 + 5 = 11
			(Addr == 'd10) ? 'b0001_000_111_000_000: // add R0 =R7 +R0 = 0
			(Addr == 'd11) ? 'b0000_010_010_100_000: // nop
			(Addr == 'd12) ? 'b0001_011_011_000_000: // add R3 =R3 +R0 = 10
			(Addr == 'd13) ? 'b0001_100_001_100_000: // add R4 =R1 +R4 = -1
			(Addr == 'd14) ? 'b0010_001_001_010_000: // SUB R1 =R1 - R2 = 10	
			(Addr == 'd15) ? 'b0011_001_001_110_000: // AND R1 =R1 &R6 = 00000010= 2
			(Addr == 'd16) ? 'b0100_001_100_001_000: // OR  R1 =R4 |R1 = 111111 = -1
			(Addr == 'd17) ? 'b0101_001_011_001_000: // XOR R1 =R3^R1 = 110101 = -11
			(Addr == 'd18) ? 'b1001_010_000_000_010: // Adi R2 = 2
			(Addr == 'd19) ? 'b0110_001_001_010_000: // SL  R1 =R1 <<R2 = 11010100
			(Addr == 'd20) ? 'b1001_010_010_000_010: // Adi R2 = R2 + 2 = 4 
			(Addr == 'd21) ? 'b1001_011_000_111_100: // Adi R3 = -4
			(Addr == 'd22) ? 'b0111_001_001_010_000: // SR  R1 =R1 >>R2 = 11111101 
			(Addr == 'd23) ? 'b1001_001_000_001_111: // addi r1 = 15
			(Addr == 'd24) ? 'b1011_011_001_111_011: // ST  Mem(R1-5 = 10) <- R3 = -4
			(Addr == 'd25) ? 'b1010_111_011_001_110: // Ld  R7 <- Mem(14 + R3 = 10) = -4
			(Addr == 'd26) ? 'b1010_110_111_001_110: // Ld  R6 <- Mem(14 + R7 = 4) = -4
			(Addr == 'd27) ? 'b0001_011_110_111_000: // Add R3 = R6 + R7 = -8
			(Addr == 'd28) ? 'b1011_011_110_000_100: // ST  Mem(R6 + 4 = 0) <- R3 = -8
			(Addr == 'd29) ? 'b1010_001_000_000_000: // Ld  R1 <- Mem(0 + R0 = 0) = -8
			(Addr == 'd30) ? 'b1001_010_000_111_011: // Adi R2 = -5
			(Addr == 'd31) ? 'b1001_001_000_000_000: // Adi R1 = 0
			(Addr == 'd32) ? 'b1100_000_001_000_001: // BR  R1 , 1 , YES
			(Addr == 'd33) ? 'b1001_010_000_000_000: // Adi R2 = 0	
			(Addr == 'd34) ? 'b1100_000_010_111_111: // BR  R2 , -1 , NOT	
			(Addr == 'd35) ? 'b1001_001_000_000_001: // Adi R1 = 1	
			(Addr == 'd36) ? 'b1100_000_001_111_011: // BR  R1 , -5 , NOT	
			(Addr == 'd37) ? 'b1100_000_000_000_000: // BR  R0 , 0 , YES	
			(Addr == 'd38) ? 'b1100_000_001_111_011: // BR  R1 , -5 , NOT 
			(Addr == 'd39) ? 'b1100_000_000_111_111: // BR  R0 , -1 , YES	
							 'b0000_000_000_000000;
					 
					 
					 /*
					 (Addr == 'd1) ? 'h1098 : //add 3, 4 -> 7
					 (Addr == 'd2) ? 'h20E0 : //sub 3, 4 -> F
					 (Addr == 'd3) ? 'h3098 : //and 3, 4 -> 0
					 (Addr == 'd4) ? 'h41D0 : //or  15, 3 -> F
					 (Addr == 'd5) ? 'h81B8 : //SRU 0x8000, 15 -> F
					 (Addr == 'd6) ? 'h71B8 : //SR 0x8000, 15 -> 1
					 */
  
  /*
  always @(*) begin
    if (set)
      //$readmemb("inst_mem.txt", InstMem);
    else
      Inst <= InstMem[Addr];
  end
  */
endmodule