module FU(
			input [2:0] id_ex_read_addr1, id_ex_read_addr2,
			ex_mem_rd, mem_wb_rd,
			input ex_mem_wb_en, mem_wb_wb_en,
			output [1:0] alu_src_sel1, alu_src_sel2);
			
			

endmodule 